VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sar_logic
  CLASS BLOCK ;
  FOREIGN sar_logic ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 246.000 73.970 250.000 ;
    END
  END clk
  PIN comp_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 246.000 77.190 250.000 ;
    END
  END comp_in
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 246.000 1.750 250.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 246.000 35.790 250.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 246.000 39.470 250.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 246.000 42.690 250.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 246.000 46.370 250.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 246.000 49.590 250.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 246.000 53.270 250.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 246.000 56.490 250.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 246.000 60.170 250.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 246.000 63.390 250.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 246.000 67.070 250.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 246.000 4.970 250.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 246.000 70.290 250.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 246.000 8.190 250.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 246.000 11.870 250.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 246.000 15.090 250.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 246.000 18.770 250.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 246.000 21.990 250.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 246.000 25.670 250.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 246.000 28.890 250.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 246.000 32.570 250.000 ;
    END
  END io_oeb[9]
  PIN output_for_analog[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END output_for_analog[0]
  PIN output_for_analog[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END output_for_analog[10]
  PIN output_for_analog[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 246.000 87.770 250.000 ;
    END
  END output_for_analog[11]
  PIN output_for_analog[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END output_for_analog[12]
  PIN output_for_analog[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 246.000 90.990 250.000 ;
    END
  END output_for_analog[13]
  PIN output_for_analog[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 246.000 94.670 250.000 ;
    END
  END output_for_analog[14]
  PIN output_for_analog[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END output_for_analog[15]
  PIN output_for_analog[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END output_for_analog[16]
  PIN output_for_analog[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 156.440 100.000 157.040 ;
    END
  END output_for_analog[17]
  PIN output_for_analog[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 219.000 100.000 219.600 ;
    END
  END output_for_analog[18]
  PIN output_for_analog[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 246.000 97.890 250.000 ;
    END
  END output_for_analog[19]
  PIN output_for_analog[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 246.000 80.870 250.000 ;
    END
  END output_for_analog[1]
  PIN output_for_analog[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END output_for_analog[2]
  PIN output_for_analog[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 246.000 84.090 250.000 ;
    END
  END output_for_analog[3]
  PIN output_for_analog[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END output_for_analog[4]
  PIN output_for_analog[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.320 100.000 31.920 ;
    END
  END output_for_analog[5]
  PIN output_for_analog[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END output_for_analog[6]
  PIN output_for_analog[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END output_for_analog[7]
  PIN output_for_analog[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 93.880 100.000 94.480 ;
    END
  END output_for_analog[8]
  PIN output_for_analog[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END output_for_analog[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.550 10.640 21.150 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.855 10.640 80.455 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 236.725 ;
      LAYER met1 ;
        RECT 1.450 10.640 97.910 236.880 ;
      LAYER met2 ;
        RECT 2.030 245.720 4.410 246.570 ;
        RECT 5.250 245.720 7.630 246.570 ;
        RECT 8.470 245.720 11.310 246.570 ;
        RECT 12.150 245.720 14.530 246.570 ;
        RECT 15.370 245.720 18.210 246.570 ;
        RECT 19.050 245.720 21.430 246.570 ;
        RECT 22.270 245.720 25.110 246.570 ;
        RECT 25.950 245.720 28.330 246.570 ;
        RECT 29.170 245.720 32.010 246.570 ;
        RECT 32.850 245.720 35.230 246.570 ;
        RECT 36.070 245.720 38.910 246.570 ;
        RECT 39.750 245.720 42.130 246.570 ;
        RECT 42.970 245.720 45.810 246.570 ;
        RECT 46.650 245.720 49.030 246.570 ;
        RECT 49.870 245.720 52.710 246.570 ;
        RECT 53.550 245.720 55.930 246.570 ;
        RECT 56.770 245.720 59.610 246.570 ;
        RECT 60.450 245.720 62.830 246.570 ;
        RECT 63.670 245.720 66.510 246.570 ;
        RECT 67.350 245.720 69.730 246.570 ;
        RECT 70.570 245.720 73.410 246.570 ;
        RECT 74.250 245.720 76.630 246.570 ;
        RECT 77.470 245.720 80.310 246.570 ;
        RECT 81.150 245.720 83.530 246.570 ;
        RECT 84.370 245.720 87.210 246.570 ;
        RECT 88.050 245.720 90.430 246.570 ;
        RECT 91.270 245.720 94.110 246.570 ;
        RECT 94.950 245.720 97.330 246.570 ;
        RECT 1.480 4.280 97.880 245.720 ;
        RECT 1.480 4.000 16.370 4.280 ;
        RECT 17.210 4.000 49.490 4.280 ;
        RECT 50.330 4.000 82.610 4.280 ;
        RECT 83.450 4.000 97.880 4.280 ;
      LAYER met3 ;
        RECT 4.000 232.920 96.000 236.805 ;
        RECT 4.400 231.520 96.000 232.920 ;
        RECT 4.000 220.000 96.000 231.520 ;
        RECT 4.000 218.600 95.600 220.000 ;
        RECT 4.000 196.880 96.000 218.600 ;
        RECT 4.400 195.480 96.000 196.880 ;
        RECT 4.000 161.520 96.000 195.480 ;
        RECT 4.400 160.120 96.000 161.520 ;
        RECT 4.000 157.440 96.000 160.120 ;
        RECT 4.000 156.040 95.600 157.440 ;
        RECT 4.000 125.480 96.000 156.040 ;
        RECT 4.400 124.080 96.000 125.480 ;
        RECT 4.000 94.880 96.000 124.080 ;
        RECT 4.000 93.480 95.600 94.880 ;
        RECT 4.000 90.120 96.000 93.480 ;
        RECT 4.400 88.720 96.000 90.120 ;
        RECT 4.000 54.080 96.000 88.720 ;
        RECT 4.400 52.680 96.000 54.080 ;
        RECT 4.000 32.320 96.000 52.680 ;
        RECT 4.000 30.920 95.600 32.320 ;
        RECT 4.000 18.720 96.000 30.920 ;
        RECT 4.400 17.320 96.000 18.720 ;
        RECT 4.000 10.715 96.000 17.320 ;
      LAYER met4 ;
        RECT 21.550 10.640 33.970 236.880 ;
        RECT 36.370 10.640 48.800 236.880 ;
        RECT 51.200 10.640 63.625 236.880 ;
        RECT 66.025 10.640 78.455 236.880 ;
        RECT 80.855 10.640 88.025 236.880 ;
  END
END sar_logic
END LIBRARY

