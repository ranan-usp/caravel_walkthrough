
module hold ( input wire comp_in,
                input wire sample,
                input wire d1b,
                input wire d2b,
                input wire d3b,
                input wire d4b,
                input wire d5b,
                input wire d6b,
                output wire r5,
                output wire r4,
                output wire r3,
                output wire r2,
                output wire r1,
                output wire r0);

    dff  dff5 ( .d(comp_in),
                .rst (sample),
                .clk (d6b),
                .q (r5),
				.qn ()),
        dff4 ( .d(comp_in),
                .rst (sample),
                .clk (d5b),
                .q (r4),
				.qn ()),
        dff3 ( .d(comp_in),
                .rst (sample),
                .clk (d4b),
                .q (r3),
				.qn ()),
        dff2 ( .d(comp_in),
                .rst (sample),
                .clk (d3b),
                .q (r2),
				.qn ()),
        dff1 ( .d(comp_in),
                .rst (sample),
                .clk (d2b),
                .q (r1),
				.qn ()),
        dff0 ( .d(comp_in),
                .rst (sample),
                .clk (d1b),
                .q (r0),
				.qn ());



endmodule